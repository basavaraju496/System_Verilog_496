`include "mcs_dv05_ADDER_Transaction.sv"
`include "mcs_dv05_ADDER_Generator.sv"
`include "mcs_dv05_ADDER_Interface.sv"
`include "mcs_dv05_ADDER_Driver.sv"
`include "mcs_dv05_ADDER_DUTMonitor.sv"
`include "mcs_dv05_ADDER_TBMonitor.sv"
`include "mcs_dv05_ADDER_Scoreboard.sv"
`include "mcs_dv05_ADDER_Coverage.sv"
`include "mcs_dv05_ADDER_Environment.sv"
`include "mcs_dv05_ADDER_Test.sv"
`include "mcs_dv05_ADDER_Top.sv"
`include "mcs_dv05_ADDER_Design.sv"
