`include"dff_dut.v"
`include"1.transaction.sv"
`include"generator.sv"
`include"interface.sv"
`include"driver.sv"
`include"ip_monitor.sv"
`include"output_monitor.sv"
`include"scoreboard.sv"
`include"environment.sv"
`include"test.sv"
`include"top.sv"
