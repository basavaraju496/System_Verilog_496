`include"1_transaction.sv"

`include"2_generator.sv"   // do var

`include"3_interface.sv"   // do var with delays

`include"4_driver.sv"   // 

`include"5_ip_monitor.sv"   // 

`include"6_dut_monitor.sv"   // 

`include"7_score_board.sv"   // 

`include "8_env.sv"

`include "test.sv"

`include "top_mux.sv"

