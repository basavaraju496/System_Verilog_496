`include "A5_Q5_Interface.sv"
`include "A5_Q5_Transaction.sv"
`include "A5_Q5_Generator.sv"
`include "A5_Q5_Driver.sv"
`include "A5_Q5_TB_monitor.sv"
`include "A5_Q5_DUT_monitor.sv"
`include "A5_Q5_Scoreboard.sv"
`include "A5_Q5_Environment.sv"
`include "A5_Q5_Test.sv"
`include "A5_Q5_top.sv"

