`include"mux8by1.v"
`include"1_transaction.sv"
`include"2_generator.sv"
`include"3_interface.sv"
`include"4_driver.sv"
`include"5_ip_monitor.sv"
`include"6_op_monitor.sv"
`include"7_score_board.sv"
`include"8_env.sv"
`include"test_mux.sv"
`include"top_mux.sv"


/*
1_transaction.sv 
3_interface.sv 
5_ip_monitor.sv 
7_score_board.sv  
Makefile 
Package.sv 
test_mux.sv 
top_mux.sv
2_generator.sv  
4_driver.sv 
6_op_monitor.sv 
8_env.sv        
mux8by1.v 
read.me  
test.sv
*/
